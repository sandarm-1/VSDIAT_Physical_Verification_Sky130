** sch_path: /home/darunix/VSDIAT_Courses/VSDIAT_PV_Sky130_3/inverter_new/xschem/inverter_new_tb.sch
**.subckt inverter_new_tb out in
*.opin out
*.opin in
x1 in net1 GND out inverter_new
V1 in GND pwl (0 0 20n 0 900n 1.8)
V2 net1 GND 1.8
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.control
tran 1n 1u
plot V(in) V(out)
.endc

**** end user architecture code
**.ends

.include inverter_new.spice
.GLOBAL GND
.end
