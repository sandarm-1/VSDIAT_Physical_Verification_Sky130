magic
tech sky130A
timestamp 1642763504
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1642674852
transform 1 0 223 0 1 -6
box -19 -24 65 296
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1642674852
transform 1 0 -7 0 1 -6
box -19 -24 249 296
<< end >>
