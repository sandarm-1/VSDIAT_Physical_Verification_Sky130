magic
tech sky130A
magscale 1 2
timestamp 1642787575
<< error_p >>
rect -52 -170 -40 -164
rect -64 -188 -62 -176
rect -64 -448 -62 -436
rect -52 -460 -40 -456
<< locali >>
rect 976 548 1936 554
rect 976 240 1622 548
rect 1930 240 1936 548
rect 976 234 1936 240
rect 334 -166 528 -142
rect -62 -176 34 -170
rect -62 -448 -52 -176
rect 20 -448 34 -176
rect 334 -322 362 -166
rect 502 -322 528 -166
rect 334 -344 528 -322
rect -62 -456 34 -448
<< viali >>
rect 1622 240 1930 548
rect -52 -448 20 -176
rect 362 -322 502 -166
rect 900 -224 968 -156
<< metal1 >>
rect 1610 548 1942 554
rect 1610 240 1622 548
rect 1930 240 1942 548
rect 1610 234 1942 240
rect 1616 -52 1936 234
rect 2222 -52 2542 -46
rect 334 -166 528 -142
rect -62 -176 34 -170
rect -62 -448 -52 -176
rect 20 -448 34 -176
rect 334 -322 362 -166
rect 502 -322 528 -166
rect 888 -156 980 -144
rect 888 -224 900 -156
rect 968 -224 980 -156
rect 888 -236 980 -224
rect 1488 -238 1558 -166
rect 334 -344 528 -322
rect 1616 -372 2222 -52
rect 2222 -378 2542 -372
rect -62 -456 34 -448
rect 1444 -570 1924 -478
rect 1832 -890 1924 -570
rect 1826 -982 1832 -890
rect 1924 -982 1930 -890
<< via1 >>
rect 2222 -372 2542 -52
rect 1832 -982 1924 -890
<< metal2 >>
rect 2222 381 2542 386
rect 2218 71 2227 381
rect 2537 71 2546 381
rect 2222 -52 2542 71
rect 2216 -372 2222 -52
rect 2542 -372 2548 -52
rect 1832 -890 1924 -884
rect 1924 -982 2432 -890
rect 1832 -988 1924 -982
rect 2340 -1142 2432 -982
rect 2760 -1142 2852 -1133
rect 2340 -1234 2760 -1142
rect 2760 -1243 2852 -1234
<< via2 >>
rect 2227 71 2537 381
rect 2760 -1234 2852 -1142
<< metal3 >>
rect 2881 386 3199 391
rect 2222 385 3200 386
rect 2222 381 2881 385
rect 2222 71 2227 381
rect 2537 71 2881 381
rect 2222 67 2881 71
rect 3199 67 3200 385
rect 2222 66 3200 67
rect 2881 61 3199 66
rect 2862 -404 2954 -398
rect 2862 -586 2954 -496
rect 2760 -678 2954 -586
rect 2760 -1137 2852 -678
rect 2755 -1142 2857 -1137
rect 2755 -1234 2760 -1142
rect 2852 -1234 2857 -1142
rect 2755 -1239 2857 -1234
<< via3 >>
rect 2881 67 3199 385
rect 2862 -496 2954 -404
<< metal4 >>
rect 2880 385 4534 386
rect 2880 67 2881 385
rect 3199 362 4534 385
rect 3199 90 4238 362
rect 4510 90 4534 362
rect 3199 67 4534 90
rect 2880 66 4534 67
rect 2861 -404 2955 -403
rect 2861 -496 2862 -404
rect 2954 -496 3190 -404
rect 2861 -497 2955 -496
<< via4 >>
rect 4238 90 4510 362
rect 3190 -610 3510 -290
<< metal5 >>
rect 4214 362 4534 386
rect 4214 90 4238 362
rect 4510 90 4534 362
rect 3166 -290 3534 -266
rect 4214 -290 4534 90
rect 3166 -610 3190 -290
rect 3510 -610 4534 -290
rect 3166 -634 3534 -610
<< labels >>
flabel space -32 16 -32 16 0 FreeSans 320 0 0 0 Exercise_2a
flabel space -14 -74 -14 -74 0 FreeSans 320 0 0 0 Via_size
flabel space 440 14 440 14 0 FreeSans 320 0 0 0 Exercise_2b
flabel space 438 -66 438 -66 0 FreeSans 320 0 0 0 Multiple_vias
flabel space 948 4 948 4 0 FreeSans 320 0 0 0 Exercise_2c
flabel space 938 -68 938 -68 0 FreeSans 320 0 0 0 Via_overlap
flabel space 1540 -4 1540 -4 0 FreeSans 320 0 0 0 Exercise_2d
flabel space 1534 -66 1534 -66 0 FreeSans 320 0 0 0 Auto_generate_via
<< end >>
