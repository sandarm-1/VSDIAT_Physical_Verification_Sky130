magic
tech sky130A
magscale 1 2
timestamp 1642789028
<< locali >>
rect -383 412 -188 446
<< viali >>
rect -417 412 -383 446
<< metal1 >>
rect 882 624 1192 698
rect 882 544 1012 624
rect 1086 544 1192 624
rect -432 455 -368 462
rect -432 403 -426 455
rect -374 403 -368 455
rect 882 442 1192 544
rect -432 396 -368 403
<< via1 >>
rect -426 446 -374 455
rect -426 412 -417 446
rect -417 412 -383 446
rect -383 412 -374 446
rect -426 403 -374 412
<< metal2 >>
rect -527 573 -383 607
rect -417 462 -383 573
rect -432 455 -368 462
rect -432 403 -426 455
rect -374 403 -368 455
rect -432 396 -368 403
<< metal4 >>
rect 16 590 146 682
<< labels >>
flabel space 70 912 70 912 0 FreeSans 320 0 0 0 Exercise_3a
flabel space 64 828 64 828 0 FreeSans 320 0 0 0 Minimum_area_rule
flabel space 1042 944 1042 944 0 FreeSans 320 0 0 0 Exercise_3b
flabel space 1018 844 1018 844 0 FreeSans 320 0 0 0 Minimum_hole_rule
flabel space 1000 334 1000 334 0 FreeSans 320 0 0 0 *must_use_drc_style_sky130(full)*
<< end >>
