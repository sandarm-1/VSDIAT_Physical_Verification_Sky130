magic
tech sky130A
magscale 1 2
timestamp 1642790788
<< dnwell >>
rect 2342 -998 3476 114
rect 5070 -1320 7036 482
<< nwell >>
rect 4990 276 7116 562
rect 2260 -124 3558 196
rect -316 -482 -26 -144
rect 640 -436 890 -178
rect 2260 -702 2642 -124
rect 3158 -702 3558 -124
rect 2260 -1080 3558 -702
rect 4990 -1114 5276 276
rect 6830 -1114 7116 276
rect 4990 -1400 7116 -1114
<< pwell >>
rect 44 -434 294 -176
rect 960 -428 1210 -170
<< psubdiff >>
rect 1112 -392 1172 -216
<< nsubdiff >>
rect 5027 505 7079 525
rect 5027 471 5107 505
rect 6999 471 7079 505
rect 5027 451 7079 471
rect 5027 445 5101 451
rect 2410 -8 2598 68
rect -260 -230 -148 -192
rect -260 -406 -228 -230
rect -176 -406 -148 -230
rect 682 -244 752 -214
rect 682 -374 698 -244
rect 738 -374 752 -244
rect 682 -400 752 -374
rect -260 -438 -148 -406
rect 2410 -898 2466 -8
rect 2540 -898 2598 -8
rect 2410 -960 2598 -898
rect 5027 -1283 5047 445
rect 5081 -1283 5101 445
rect 5027 -1289 5101 -1283
rect 7005 445 7079 451
rect 7005 -1283 7025 445
rect 7059 -1283 7079 445
rect 7005 -1289 7079 -1283
rect 5027 -1309 7079 -1289
rect 5027 -1343 5107 -1309
rect 6999 -1343 7079 -1309
rect 5027 -1363 7079 -1343
<< nsubdiffcont >>
rect 5107 471 6999 505
rect -228 -406 -176 -230
rect 698 -374 738 -244
rect 2466 -898 2540 -8
rect 5047 -1283 5081 445
rect 7025 -1283 7059 445
rect 5107 -1343 6999 -1309
<< locali >>
rect 5047 471 5107 505
rect 6999 471 7059 505
rect 5047 445 5081 471
rect 2460 -8 2544 22
rect -234 -230 -172 -212
rect -234 -406 -228 -230
rect -176 -406 -172 -230
rect 682 -244 752 -214
rect 682 -374 698 -244
rect 738 -374 752 -244
rect 682 -400 752 -374
rect -234 -432 -172 -406
rect 2460 -898 2466 -8
rect 2540 -898 2544 -8
rect 2460 -938 2544 -898
rect 5047 -1309 5081 -1283
rect 7025 445 7059 471
rect 7025 -1309 7059 -1283
rect 5047 -1343 5107 -1309
rect 6999 -1343 7059 -1309
<< labels >>
flabel space -28 8 -28 8 0 FreeSans 320 0 0 0 Exercise_4a
flabel space -26 -68 -26 -68 0 FreeSans 320 0 0 0 Wells
flabel space 926 -16 926 -16 0 FreeSans 320 0 0 0 Exercise_4b
flabel space 920 -84 920 -84 0 FreeSans 320 0 0 0 Wells
flabel space 1936 68 1936 68 0 FreeSans 320 0 0 0 Exercise_4c
flabel space 1922 -8 1922 -8 0 FreeSans 320 0 0 0 Deep_NWell
<< end >>
